module Add_FSM(
    input clock,
    input reset,
    output done
)


