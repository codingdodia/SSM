module Add_FSM(
    input clock,
    input reset,
    input [6:0] param1;
    input [6:0] param2;
    output done
);




